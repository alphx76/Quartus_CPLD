-- DI seno e
compuerta or
library IEEE;
_ LOGIC_1164. ALL ;
use IEEE.STD
use IEEE.
use
aentity proyectol is
a port (A
B
x
end entity;
. in STD_LOGIC;
. in STD_LOG1q,•
. out STD_LOGIC);
aarchitecture compuerta_or of proyectol is
abegin
salida<= entradal
entrada2;
or
end architecture;